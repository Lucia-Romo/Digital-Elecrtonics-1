----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:37:34 04/30/2020 
-- Design Name: 
-- Module Name:    binary_cnt - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;    -- Provides unsigned numerical computation

------------------------------------------------------------------------
-- Entity declaration for N-bit binary counter
------------------------------------------------------------------------
entity binary_cnt is
generic (
    g_NBIT : positive := 4      -- Number of bits
);
port (
    clk_i     : in  std_logic;
    srst_n_i  : in  std_logic;   -- Synchronous reset (active low)
    en_i      : in  std_logic;   -- Enable
	 in_encoder:in  std_logic_vector(g_NBIT-1 downto 0);
	 
    cnt_o     : out std_logic_vector(g_NBIT-1 downto 0)
);
end entity binary_cnt;

architecture Behavioral of binary_cnt is

	signal s_cnt : std_logic_vector(g_NBIT-1 downto 0);

	begin
	   
	s_cnt <= in_encoder;
	
    --------------------------------------------------------------------
    -- p_binary_cnt:
    -- Sequential process with synchronous reset and clock enable,
    -- which implements a one-way binary counter.
    --------------------------------------------------------------------
    p_binary_cnt : process (clk_i, en_i)

    begin
        if rising_edge(clk_i) then  -- Rising clock edge
            if srst_n_i = '0' then  -- Synchronous reset (active low)
                s_cnt <= (others => '1');   --Initialization at "1111"
					 elsif en_i = '1' then
                s_cnt <= s_cnt - 1; -- Normal operation
            end if;
        end if;
    end process p_binary_cnt;

    cnt_o <= s_cnt;

		

end Behavioral;

